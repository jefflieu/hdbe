
`define OPCODE_ADD    "     add"
`define OPCODE_SUB    "     sub"
`define OPCODE_OR     "      or"
`define OPCODE_AND    "     and"
`define OPCODE_XOR    "     xor"
`define OPCODE_MUL    "     mul"
`define OPCODE_ADD    "     add"
`define OPCODE_LSHR   "    lshr"
`define OPCODE_ASHR   "    ashr"
`define OPCODE_SHL    "     shl"
`define OPCODE_ZEXT   "    zext"
`define OPCODE_SEXT   "    sext"
`define OPCODE_TRUNC  "   trunc"
`define OPCODE_EQ     "      eq"
`define OPCODE_NE     "      ne"
`define OPCODE_UGT    "     ugt"
`define OPCODE_ULT    "     ult"
`define OPCODE_UGE    "     uge"
`define OPCODE_ULE    "     ule"
`define OPCODE_SGT    "     ugt"
`define OPCODE_SLT    "     ult"
`define OPCODE_SGE    "     uge"
`define OPCODE_SLE    "     ule"
